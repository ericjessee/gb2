`define TEST_MEM_DEPTH 16'h3f46 //gameboy rom size
`define PC_INIT 16'h0001
`define SP_INIT `TEST_MEM_DEPTH