typedef enum logic [7:0] {
    OP_NOP          = 8'h00,
    OP_LD_BC_D16    = 8'h01,
    OP_LDPTR_BC_A   = 8'h02,
    OP_INC_BC       = 8'h03,
    OP_INC_B        = 8'h04,
    OP_DEC_B        = 8'h05,
    OP_LD_B_D8      = 8'h06,
    OP_RLCA         = 8'h07,
    OP_LDPTR_A16_SP = 8'h08,
    OP_ADD_HL_BC    = 8'h09,
    OP_LDPTR_A_BC   = 8'h0a,
    OP_DEC_BC       = 8'h0b,
    OP_INC_C        = 8'h0c,
    OP_DEC_C        = 8'h0d,
    OP_LD_C_D8      = 8'h0e,
    OP_RRCA         = 8'h0f,
    OP_STOP         = 8'h10,
    OP_LD_DE_D16    = 8'h11,
    OP_LDPTR_DE_A   = 8'h12,
    OP_INC_DE       = 8'h13,
    OP_INC_D        = 8'h14,
    OP_DEC_D        = 8'h15,
    OP_LD_D_D8      = 8'h16,
    OP_RLA          = 8'h17,
    OP_JR_S8        = 8'h18,
    OP_ADD_HL_DE    = 8'h19,
    OP_LDPTR_A_DE   = 8'h1a,
    OP_DEC_DE       = 8'h1b,
    OP_INC_E        = 8'h1c,
    OP_DEC_E        = 8'h1d,
    OP_LD_E_D8      = 8'h1e,
    OP_RRA          = 8'h1f,
    OP_JR_NZ_S8     = 8'h20,
    OP_LD_HL_D16    = 8'h21,
    OP_LDPTR_HLI_A  = 8'h22,
    OP_INC_HL       = 8'h23,
    OP_INC_H        = 8'h24,
    OP_DEC_H        = 8'h25,
    OP_LD_H_D8      = 8'h26,
    OP_DAA          = 8'h27,
    OP_JR_Z_S8      = 8'h28,
    OP_ADD_HL_HL    = 8'h29,
    OP_LDPTR_A_HLI  = 8'h2a,
    OP_DEC_HL       = 8'h2b,
    OP_INC_L        = 8'h2c,
    OP_DEC_L        = 8'h2d,
    OP_LD_L_D8      = 8'h2e,
    OP_CPL          = 8'h2f,
    OP_JR_NC_S8     = 8'h30,
    OP_LD_SP_D16    = 8'h31,
    OP_LDPTR_HLD_A  = 8'h32,
    OP_INC_SP       = 8'h33,
    OP_INCPTR_HL    = 8'h34,
    OP_DECPTR_HL    = 8'h35,
    OP_LDPTR_HL_D8  = 8'h36,
    OP_SCF          = 8'h37,
    OP_JR_C_S8      = 8'h38,
    OP_ADD_HL_SP    = 8'h39,
    OP_LDPTR_A_HLD  = 8'h3a,
    OP_DEC_SP       = 8'h3b,
    OP_INC_A        = 8'h3c,
    OP_DEC_A        = 8'h3d,
    OP_LD_A_D8      = 8'h3e,
    OP_CCF          = 8'h3f,
    OP_LD_B_B       = 8'h40,
    OP_LD_B_C       = 8'h41,
    OP_LD_B_D       = 8'h42,
    OP_LD_B_E       = 8'h43,
    OP_LD_B_H       = 8'h44,
    OP_LD_B_L       = 8'h45,
    OP_LDPTR_B_HL   = 8'h46,
    OP_LD_B_A       = 8'h47,
    OP_LD_C_B       = 8'h48,
    OP_LD_C_C       = 8'h49,
    OP_LD_C_D       = 8'h4a,
    OP_LD_C_E       = 8'h4b,
    OP_LD_C_H       = 8'h4c,
    OP_LD_C_L       = 8'h4d,
    OP_LDPTR_C_HL   = 8'h4e,
    OP_LD_C_A       = 8'h4f,
    OP_LD_D_B       = 8'h50,
    OP_LD_D_C       = 8'h51,
    OP_LD_D_D       = 8'h52,
    OP_LD_D_E       = 8'h53,
    OP_LD_D_H       = 8'h54,
    OP_LD_D_L       = 8'h55,
    OP_LDPTR_D_HL   = 8'h56,
    OP_LD_D_A       = 8'h57,
    OP_LD_E_B       = 8'h58,
    OP_LD_E_C       = 8'h59,
    OP_LD_E_D       = 8'h5a,
    OP_LD_E_E       = 8'h5b,
    OP_LD_E_H       = 8'h5c,
    OP_LD_E_L       = 8'h5d,
    OP_LDPTR_E_HL   = 8'h5e,
    OP_LD_E_A       = 8'h5f,
    OP_LD_H_B       = 8'h60,
    OP_LD_H_C       = 8'h61,
    OP_LD_H_D       = 8'h62,
    OP_LD_H_E       = 8'h63,
    OP_LD_H_H       = 8'h64,
    OP_LD_H_L       = 8'h65,
    OP_LDPTR_H_HL   = 8'h66,
    OP_LD_H_A       = 8'h67,
    OP_LD_L_B       = 8'h68,
    OP_LD_L_C       = 8'h69,
    OP_LD_L_D       = 8'h6a,
    OP_LD_L_E       = 8'h6b,
    OP_LD_L_H       = 8'h6c,
    OP_LD_L_L       = 8'h6d,
    OP_LDPTR_L_HL   = 8'h6e,
    OP_LD_L_A       = 8'h6f,
    OP_LDPTR_HL_B   = 8'h70,
    OP_LDPTR_HL_C   = 8'h71,
    OP_LDPTR_HL_D   = 8'h72,
    OP_LDPTR_HL_E   = 8'h73,
    OP_LDPTR_HL_H   = 8'h74,
    OP_LDPTR_HL_L   = 8'h75,
    OP_HALT         = 8'h76,
    OP_LDPTR_HL_A   = 8'h77,
    OP_LD_A_B       = 8'h78,
    OP_LD_A_C       = 8'h79,
    OP_LD_A_D       = 8'h7a,
    OP_LD_A_E       = 8'h7b,
    OP_LD_A_H       = 8'h7c,
    OP_LD_A_L       = 8'h7d,
    OP_LDPTR_A_HL   = 8'h7e,
    OP_LD_A_A       = 8'h7f,
    OP_ADD_A_B      = 8'h80,
    OP_ADD_A_C      = 8'h81,
    OP_ADD_A_D      = 8'h82,
    OP_ADD_A_E      = 8'h83,
    OP_ADD_A_H      = 8'h84,
    OP_ADD_A_L      = 8'h85,
    OP_ADDPTR_A_HL  = 8'h86,
    OP_ADD_A_A      = 8'h87,
    OP_ADC_A_B      = 8'h88,
    OP_ADC_A_C      = 8'h89,
    OP_ADC_A_D      = 8'h8a,
    OP_ADC_A_E      = 8'h8b,
    OP_ADC_A_H      = 8'h8c,
    OP_ADC_A_L      = 8'h8d,
    OP_ADCPTR_A_HL  = 8'h8e,
    OP_ADC_A_A      = 8'h8f,
    OP_SUB_A_B      = 8'h90,
    OP_SUB_A_C      = 8'h91,
    OP_SUB_A_D      = 8'h92,
    OP_SUB_A_E      = 8'h93,
    OP_SUB_A_H      = 8'h94,
    OP_SUB_A_L      = 8'h95,
    OP_SUBPTR_A_HL  = 8'h96,
    OP_SUB_A_A      = 8'h97,
    OP_SBC_A_B      = 8'h98,
    OP_SBC_A_C      = 8'h99,
    OP_SBC_A_D      = 8'h9a,
    OP_SBC_A_E      = 8'h9b,
    OP_SBC_A_H      = 8'h9c,
    OP_SBC_A_L      = 8'h9d,
    OP_SBCPTR_A_HL  = 8'h9e,
    OP_SBC_A_A      = 8'h9f,
    OP_AND_A_B      = 8'ha0,
    OP_AND_A_C      = 8'ha1,
    OP_AND_A_D      = 8'ha2,
    OP_AND_A_E      = 8'ha3,
    OP_AND_A_H      = 8'ha4,
    OP_AND_A_L      = 8'ha5,
    OP_ANDPTR_A_HL  = 8'ha6,
    OP_AND_A_A      = 8'ha7,
    OP_XOR_A_B      = 8'ha8,
    OP_XOR_A_C      = 8'ha9,
    OP_XOR_A_D      = 8'haa,
    OP_XOR_A_E      = 8'hab,
    OP_XOR_A_H      = 8'hac,
    OP_XOR_A_L      = 8'had,
    OP_XORPTR_A_HL  = 8'hae,
    OP_XOR_A_A      = 8'haf,
    OP_OR_A_B       = 8'hb0,
    OP_OR_A_C       = 8'hb1,
    OP_OR_A_D       = 8'hb2,
    OP_OR_A_E       = 8'hb3,
    OP_OR_A_H       = 8'hb4,
    OP_OR_A_L       = 8'hb5,
    OP_ORPTR_A_HL   = 8'hb6,
    OP_OR_A_A       = 8'hb7,
    OP_CP_A_B       = 8'hb8,
    OP_CP_A_C       = 8'hb9,
    OP_CP_A_D       = 8'hba,
    OP_CP_A_E       = 8'hbb,
    OP_CP_A_H       = 8'hbc,
    OP_CP_A_L       = 8'hbd,
    OP_CPPTR_A_HL   = 8'hbe,
    OP_CP_A_A       = 8'hbf,
    OP_RET_NZ       = 8'hc0,
    OP_POP_BC       = 8'hc1,
    OP_JP_NZ_A16    = 8'hc2,
    OP_JP_A16       = 8'hc3,
    OP_CALL_NZ_A16  = 8'hc4,
    OP_PUSH_BC      = 8'hc5,
    OP_ADD_A_D8     = 8'hc6,
    OP_RST_0        = 8'hc7,
    OP_RET_Z        = 8'hc8,
    OP_RET          = 8'hc9,
    OP_JP_NZ_A16    = 8'hca,
    OP_INSTR_16     = 8'hcb,
    OP_CALL_Z_A16   = 8'hcc,
    OP_CALL_A16     = 8'hcd,
    OP_ADC_A_D8     = 8'hce,
    OP_RST_1        = 8'hcf,
    OP_RET_NC       = 8'hd0,
    OP_POP_DE       = 8'hd1,
    OP_JP_NC_A16    = 8'hd2,
    NULL1           = 8'hd3,
    OP_CALL_NC_A16  = 8'hd4,
    OP_PUSH_DE      = 8'hd5,
    OP_SUB_A_D8     = 8'hd6,
    OP_RST_2        = 8'hd7,
    OP_RET_C        = 8'hd8,
    OP_RETI         = 8'hd9,
    OP_JP_C_A16     = 8'hda,
    NULL2           = 8'hdb,
    OP_CALL_C_A16   = 8'hdc,
    NULL3           = 8'hdd,
    OP_SBC_A_D8     = 8'hde,
    OP_RST_3        = 8'hdf,
    OP_LDPTR_A8_A   = 8'he0,
    OP_POP_HL       = 8'he1,
    OP_LDPTR_C_A    = 8'he2,
    NULL4           = 8'he3,
    NULL5           = 8'he4,
    OP_PUSH_HL      = 8'he5,
    OP_AND_A_D8     = 8'he6,
    OP_RST_4        = 8'he7,
    OP_ADD_SP       = 8'he8,
    OP_JP_HL        = 8'he9,
    OP_LDPTR_A16_A  = 8'hea,
    NULL6           = 8'heb,
    NULL7           = 8'hec,
    NULL8           = 8'hed,
    OP_XOR_A_D8     = 8'hee,
    OP_RST_5        = 8'hef,
    OP_LDPTR_A_A8   = 8'hf0,
    OP_POP_AF       = 8'hf1,
    OP_LDPTR_A_C    = 8'hf2,
    DI              = 8'hf3,
    NULL9           = 8'hf4,
    OP_PUSH_AF      = 8'hf5,
    OP_OR_A_D8      = 8'hf6,
    OP_RST_6        = 8'hf7,
    OP_LD_HL_SP_S8  = 8'hf8,
    OP_SP_HL        = 8'hf9,
    OP_LDPTR_A_A16  = 8'hfa,
    EI              = 8'hfb,
    NULL10          = 8'hfc,
    NULL11          = 8'hfd,
    OP_CP_A_D8      = 8'hfe,
    OP_RST_7        = 8'hff
} opcode8_t;

typedef enum logic [7:0] {
    OP_RLC_B        = 8'h00,
    OP_RLC_C        = 8'h01,
    OP_RLC_D        = 8'h02,
    OP_RLC_E        = 8'h03,
    OP_RLC_H        = 8'h04,
    OP_RLC_L        = 8'h05,
    OP_RLCPTR_HL    = 8'h06,
    OP_RLC_A        = 8'h07,
    OP_RRC_B        = 8'h08,
    OP_RRC_C        = 8'h09,
    OP_RRC_D        = 8'h0a,
    OP_RRC_E        = 8'h0b,
    OP_RRC_H        = 8'h0c,
    OP_RRC_L        = 8'h0d,
    OP_RRCPTR_HL    = 8'h0e,
    OP_RRC_A        = 8'h0f,
    OP_RL_B         = 8'h10,
    OP_RL_C         = 8'h11,
    OP_RL_D         = 8'h12,
    OP_RL_E         = 8'h13,
    OP_RL_H         = 8'h14,
    OP_RL_L         = 8'h15,
    OP_RLPTR_HL     = 8'h16,
    OP_RL_A         = 8'h17,
    OP_RR_B         = 8'h18,
    OP_RR_C         = 8'h19,
    OP_RR_D         = 8'h1a,
    OP_RR_E         = 8'h1b,
    OP_RR_H         = 8'h1c,
    OP_RR_L         = 8'h1d,
    OP_RRPTR_HL     = 8'h1e,
    OP_RR_A         = 8'h1f,
    OP_SLA_B        = 8'h20,
    OP_SLA_C        = 8'h21,
    OP_SLA_D        = 8'h22,
    OP_SLA_E        = 8'h23,
    OP_SLA_H        = 8'h24,
    OP_SLA_L        = 8'h25,
    OP_SLAPTR_HL    = 8'h26,
    OP_SLA_A        = 8'h27,
    OP_SRA_B        = 8'h28,
    OP_SRA_C        = 8'h29,
    OP_SRA_D        = 8'h2a,
    OP_SRA_E        = 8'h2b,
    OP_SRA_H        = 8'h2c,
    OP_SRA_L        = 8'h2d,
    OP_SRAPTR_HL    = 8'h2e,
    OP_SRA_A        = 8'h2f,
    OP_SWAP_B       = 8'h30,
    OP_SWAP_C       = 8'h31,
    OP_SWAP_D       = 8'h32,
    OP_SWAP_E       = 8'h33,
    OP_SWAP_H       = 8'h34,
    OP_SWAP_L       = 8'h35,
    OP_SWAPPTR_HL   = 8'h36,
    OP_SWAP_A       = 8'h37,
    OP_SRL_B        = 8'h38,
    OP_SRL_C        = 8'h39,
    OP_SRL_D        = 8'h3a,
    OP_SRL_E        = 8'h3b,
    OP_SRL_H        = 8'h3c,
    OP_SRL_L        = 8'h3d,
    OP_SRLPTR_HL    = 8'h3e,
    OP_SRL_A        = 8'h3f,
    OP_BIT0_B       = 8'h40,
    OP_BIT0_C       = 8'h41,
    OP_BIT0_D       = 8'h42,
    OP_BIT0_E       = 8'h43,
    OP_BIT0_H       = 8'h44,
    OP_BIT0_L       = 8'h45,
    OP_BIT0PTR_HL   = 8'h46,
    OP_BIT0_A       = 8'h47,
    OP_BIT1_B       = 8'h48,
    OP_BIT1_C       = 8'h49,
    OP_BIT1_D       = 8'h4a,
    OP_BIT1_E       = 8'h4b,
    OP_BIT1_H       = 8'h4c,
    OP_BIT1_L       = 8'h4d,
    OP_BIT1PTR_HL   = 8'h4e,
    OP_BIT1_A       = 8'h4f,
    OP_BIT2_B       = 8'h50,
    OP_BIT2_C       = 8'h51,
    OP_BIT2_D       = 8'h52,
    OP_BIT2_E       = 8'h53,
    OP_BIT2_H       = 8'h54,
    OP_BIT2_L       = 8'h55,
    OP_BIT2PTR_HL   = 8'h56,
    OP_BIT2_A       = 8'h57,
    OP_BIT3_B       = 8'h58,
    OP_BIT3_C       = 8'h59,
    OP_BIT3_D       = 8'h5a,
    OP_BIT3_E       = 8'h5b,
    OP_BIT3_H       = 8'h5c,
    OP_BIT3_L       = 8'h5d,
    OP_BIT3PTR_HL   = 8'h5e,
    OP_BIT3_A       = 8'h5f,
    OP_BIT4_B       = 8'h60,
    OP_BIT4_C       = 8'h61,
    OP_BIT4_D       = 8'h62,
    OP_BIT4_E       = 8'h63,
    OP_BIT4_H       = 8'h64,
    OP_BIT4_L       = 8'h65,
    OP_BIT4PTR_HL   = 8'h66,
    OP_BIT4_A       = 8'h67,
    OP_BIT5_B       = 8'h68,
    OP_BIT5_C       = 8'h69,
    OP_BIT5_D       = 8'h6a,
    OP_BIT5_E       = 8'h6b,
    OP_BIT5_H       = 8'h6c,
    OP_BIT5_L       = 8'h6d,
    OP_BIT5PTR_HL   = 8'h6e,
    OP_BIT5_A       = 8'h6f,
    OP_BIT6_B       = 8'h70,
    OP_BIT6_C       = 8'h71,
    OP_BIT6_D       = 8'h72,
    OP_BIT6_E       = 8'h73,
    OP_BIT6_H       = 8'h74,
    OP_BIT6_L       = 8'h75,
    OP_BIT6PTR_HL   = 8'h76,
    OP_BIT6_A       = 8'h77,
    OP_BIT7_B       = 8'h78,
    OP_BIT7_C       = 8'h79,
    OP_BIT7_D       = 8'h7a,
    OP_BIT7_E       = 8'h7b,
    OP_BIT7_H       = 8'h7c,
    OP_BIT7_L       = 8'h7d,
    OP_BIT7PTR_HL   = 8'h7e,
    OP_BIT7_A       = 8'h7f,
    OP_RES0_B       = 8'h80,
    OP_RES0_C       = 8'h81,
    OP_RES0_D       = 8'h82,
    OP_RES0_E       = 8'h83,
    OP_RES0_H       = 8'h84,
    OP_RES0_L       = 8'h85,
    OP_RES0PTR_HL   = 8'h86,
    OP_RES0_A       = 8'h87,
    OP_RES1_B       = 8'h88,
    OP_RES1_C       = 8'h89,
    OP_RES1_D       = 8'h8a,
    OP_RES1_E       = 8'h8b,
    OP_RES1_H       = 8'h8c,
    OP_RES1_L       = 8'h8d,
    OP_RES1PTR_HL   = 8'h8e,
    OP_RES1_A       = 8'h8f,
    OP_RES2_B       = 8'h90,
    OP_RES2_C       = 8'h91,
    OP_RES2_D       = 8'h92,
    OP_RES2_E       = 8'h93,
    OP_RES2_H       = 8'h94,
    OP_RES2_L       = 8'h95,
    OP_RES2PTR_HL   = 8'h96,
    OP_RES2_A       = 8'h97,
    OP_RES3_B       = 8'h98,
    OP_RES3_C       = 8'h99,
    OP_RES3_D       = 8'h9a,
    OP_RES3_E       = 8'h9b,
    OP_RES3_H       = 8'h9c,
    OP_RES3_L       = 8'h9d,
    OP_RES3PTR_HL   = 8'h9e,
    OP_RES3_A       = 8'h9f,
    OP_RES4_B       = 8'ha0,
    OP_RES4_C       = 8'ha1,
    OP_RES4_D       = 8'ha2,
    OP_RES4_E       = 8'ha3,
    OP_RES4_H       = 8'ha4,
    OP_RES4_L       = 8'ha5,
    OP_RES4PTR_HL   = 8'ha6,
    OP_RES4_A       = 8'ha7,
    OP_RES5_B       = 8'ha8,
    OP_RES5_C       = 8'ha9,
    OP_RES5_D       = 8'haa,
    OP_RES5_E       = 8'hab,
    OP_RES5_H       = 8'hac,
    OP_RES5_L       = 8'had,
    OP_RES5PTR_HL   = 8'hae,
    OP_RES5_A       = 8'haf,
    OP_RES6_B       = 8'hb0,
    OP_RES6_C       = 8'hb1,
    OP_RES6_D       = 8'hb2,
    OP_RES6_E       = 8'hb3,
    OP_RES6_H       = 8'hb4,
    OP_RES6_L       = 8'hb5,
    OP_RES6PTR_HL   = 8'hb6,
    OP_RES6_A       = 8'hb7,
    OP_RES7_B       = 8'hb8,
    OP_RES7_C       = 8'hb9,
    OP_RES7_D       = 8'hba,
    OP_RES7_E       = 8'hbb,
    OP_RES7_H       = 8'hbc,
    OP_RES7_L       = 8'hbd,
    OP_RES7PTR_HL   = 8'hbe,
    OP_RES7_A       = 8'hbf,
    OP_SET0_B       = 8'hc0,
    OP_SET0_C       = 8'hc1,
    OP_SET0_D       = 8'hc2,
    OP_SET0_E       = 8'hc3,
    OP_SET0_H       = 8'hc4,
    OP_SET0_L       = 8'hc5,
    OP_SET0PTR_HL   = 8'hc6,
    OP_SET0_A       = 8'hc7,
    OP_SET1_B       = 8'hc8,
    OP_SET1_C       = 8'hc9,
    OP_SET1_D       = 8'hca,
    OP_SET1_E       = 8'hcb,
    OP_SET1_H       = 8'hcc,
    OP_SET1_L       = 8'hcd,
    OP_SET1PTR_HL   = 8'hce,
    OP_SET1_A       = 8'hcf,
    OP_SET2_B       = 8'hd0,
    OP_SET2_C       = 8'hd1,
    OP_SET2_D       = 8'hd2,
    OP_SET2_E       = 8'hd3,
    OP_SET2_H       = 8'hd4,
    OP_SET2_L       = 8'hd5,
    OP_SET2PTR_HL   = 8'hd6,
    OP_SET2_A       = 8'hd7,
    OP_SET3_B       = 8'hd8,
    OP_SET3_C       = 8'hd9,
    OP_SET3_D       = 8'hda,
    OP_SET3_E       = 8'hdb,
    OP_SET3_H       = 8'hdc,
    OP_SET3_L       = 8'hdd,
    OP_SET3PTR_HL   = 8'hde,
    OP_SET3_A       = 8'hdf,
    OP_SET4_B       = 8'he0,
    OP_SET4_C       = 8'he1,
    OP_SET4_D       = 8'he2,
    OP_SET4_E       = 8'he3,
    OP_SET4_H       = 8'he4,
    OP_SET4_L       = 8'he5,
    OP_SET4PTR_HL   = 8'he6,
    OP_SET4_A       = 8'he7,
    OP_SET5_B       = 8'he8,
    OP_SET5_C       = 8'he9,
    OP_SET5_D       = 8'hea,
    OP_SET5_E       = 8'heb,
    OP_SET5_H       = 8'hec,
    OP_SET5_L       = 8'hed,
    OP_SET5PTR_HL   = 8'hee,
    OP_SET5_A       = 8'hef,
    OP_SET6_B       = 8'hf0,
    OP_SET6_C       = 8'hf1,
    OP_SET6_D       = 8'hf2,
    OP_SET6_E       = 8'hf3,
    OP_SET6_H       = 8'hf4,
    OP_SET6_L       = 8'hf5,
    OP_SET6PTR_HL   = 8'hf6,
    OP_SET6_A       = 8'hf7,
    OP_SET7_B       = 8'hf8,
    OP_SET7_C       = 8'hf9,
    OP_SET7_D       = 8'hfa,
    OP_SET7_E       = 8'hfb,
    OP_SET7_H       = 8'hfc,
    OP_SET7_L       = 8'hfd,
    OP_SET7PTR_HL   = 8'hfe,
    OP_SET7_A       = 8'hff
} opcode16_t;