`define TEST_MEM_DEPTH 16'd256
`define PC_INIT 16'h0001
`define SP_INIT `TEST_MEM_DEPTH