`define TEST_MEM_DEPTH 16'hffff
`define PC_INIT 16'h0001
`define SP_INIT `TEST_MEM_DEPTH