`ifndef __GLOBAL_DEFINES_VH__
`define __GLOBAL_DEFINES_VH__

`define TEST_MEM_DEPTH 16'hffff
`define PC_INIT 16'h0000
`define SP_INIT 16'hc100

`endif
