module fetch (
    

);

endmodule